//========================================================================== //
// Copyright (c) 2022, Stephen Henry
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// * Redistributions of source code must retain the above copyright notice, this
//   list of conditions and the following disclaimer.
//
// * Redistributions in binary form must reproduce the above copyright notice,
//   this list of conditions and the following disclaimer in the documentation
//   and/or other materials provided with the distribution.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//========================================================================== //

`include "common_defs.vh"

`include "q_pkg.vh"
`include "cfg_pkg.vh"
//`include "eng/eng_pipe_xa_rom_pkg.vh"

module eng_pipe_xa (
// -------------------------------------------------------------------------- //
//
//  input eng_pipe_xa_rom_pkg::rom_pc_t             i_fa_pc_r

// -------------------------------------------------------------------------- //
// Clk/Reset
  input wire logic                                clk
, input wire logic                                arst_n
);

// ========================================================================== //
//                                                                            //
//  Instances                                                                 //
//                                                                            //
// ========================================================================== //
/*
// -------------------------------------------------------------------------- //
//
case (cfg_pkg::UCODE_TYPE)
cfg_pkg::UCODE_HOR: begin : ucode_hor_GEN

eng_pipe_xa_rom u_eng_pipe_xa_rom (
//
  .i_pc                      (i_fa_pc_r)
//
, .o_inst                    ()
);

end : ucode_hor_GEN
cfg_pkg::UCODE_VER: begin : ucode_ver_GEN

eng_pipe_xa_rom u_eng_pipe_xa_rom (
//
  .i_pc                      ()
//
, .o_inst                    ()
);

eng_pipe_xa_dec u_eng_pipe_xa_dec (
);

end : ucode_ver_GEN
endcase
*/
endmodule : eng_pipe_xa
